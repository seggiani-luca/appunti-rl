// un adder a 4 cifre in base 2 che calcola @x3_x0 + @y3_y0, 
// mettendo il risultato in @s3_s0 e il riporto in @cout, aggiornato
// con un flag di overflow @ow
module n4_b2_adder_i(x3_x0, y3_y0, cin, s3_s0, cout, ow);
	input[3:0] x3_x0, y3_y0;
	input cin;	
	output[3:0] s3_s0;
	output cout, ow;

	wire[3:0] carry;
	assign cout = carry[3];

	assign ow = carry[3] ^ carry[2];

	b2_adder add_0 (
		.x(x3_x0[0]), .y(y3_y0[0]),
		.cin(cin),
		.s(s3_s0[0]),
		.cout(carry[0])
	);
	
	b2_adder add_1 (
		.x(x3_x0[1]), .y(y3_y0[1]),
		.cin(carry[0]),
		.s(s3_s0[1]),
		.cout(carry[1])
	);

	b2_adder add_2 (
		.x(x3_x0[2]), .y(y3_y0[2]),
		.cin(carry[1]),
		.s(s3_s0[2]),
		.cout(carry[2])
	);
	
	b2_adder add_3 (
		.x(x3_x0[3]), .y(y3_y0[3]),
		.cin(carry[2]),
		.s(s3_s0[3]),
		.cout(carry[3])
	);
endmodule
