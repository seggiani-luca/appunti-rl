// un estensore di campo per interi in codifica binaria con LSD @x,
// che mette in @x_est la nuova LSD
module b2_field_extensor(x, x_est);
	input x;
	output x_est;

	assign x = x_est;
endmodule
